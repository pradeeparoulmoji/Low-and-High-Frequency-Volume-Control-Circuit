* C:\Users\prada\Desktop\PROGETTO ELETTRONICA\FINALL2 transient test.sch

* Schematics Version 9.1 - Web Update 1
* Wed Jan 10 17:54:12 2024



** Analysis setup **
.tran 0ns 1000000ns
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "FINALL2 transient test.net"
.INC "FINALL2 transient test.als"


.probe


.END
